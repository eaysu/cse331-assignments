module not32(out, a);

input [31:0] a;
output [31:0] out;

   // 32 bit not operation
	not(out[0], a[0]);
	not(out[1], a[1]);
	not(out[2], a[2]);
	not(out[3], a[3]);
	not(out[4], a[4]);
	not(out[5], a[5]);
	not(out[6], a[6]);
	not(out[7], a[7]);
	not(out[8], a[8]);
	not(out[9], a[9]);
	not(out[10], a[10]);
	not(out[11], a[11]);
	not(out[12], a[12]);
	not(out[13], a[13]);
	not(out[14], a[14]);
	not(out[15], a[15]);
	not(out[16], a[16]);
	not(out[17], a[17]);
	not(out[18], a[18]);
	not(out[19], a[19]);
	not(out[20], a[20]);
	not(out[21], a[21]);
	not(out[22], a[22]);
	not(out[23], a[23]);
	not(out[24], a[24]);
	not(out[25], a[25]);
	not(out[26], a[26]);
	not(out[27], a[27]);
	not(out[28], a[28]);
	not(out[29], a[29]);
	not(out[30], a[30]);
	not(out[31], a[31]);

endmodule