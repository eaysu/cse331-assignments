module instr_mem        
(  
      input         [15:0]     pc,  
      output wire   [31:0]     instruction  
); 
			  
      reg [31:0] rom[1023:0];  
      initial  
      begin  
	       rom[0] = 32'b01100000000001000000000000001100; // li $1, 3
          rom[1] = 32'b00000000000001000100000000000000;
          rom[2] = 32'b01100000000010000000000000010100; // li $2, 5
          rom[3] = 32'b00000000000010001000000000000000;
			 rom[4] = 32'b00000000100001010000001000100000; // sub $4, $2, $1
          rom[5] = 32'b00000000000100010000000000000000;
          rom[6] = 32'b00000000010010001100001000000000; // add $3, $2, $1
          rom[7] = 32'b00000000000011001100000000000000;
          rom[8] = 32'b01100000001000000000000000101100; // li $8, 11
          rom[9] = 32'b00000000001000100000000000000000;
			 rom[10] = 32'b01100000000111000000000000000000; // li $7, 0
          rom[11] = 32'b00000000000111011100000000000000;
          rom[12] = 32'b00100010001000111111111111111100; // addi $8, $8, -1
          rom[13] = 32'b00000000001000100011110000000000;
			 rom[14] = 32'b10101100000100000000001100100000; // sw $4, 100($0)
          rom[15] = 32'b00000000000100010000000000000000;
          rom[16] = 32'b10001100000110000000001100100000; // lw $6, 100($0)
          rom[17] = 32'b00000000000110011000000000000000;
          rom[18] = 32'b00000011100000000000000010000000; // jr $14
          rom[19] = 32'b00000000000000000000000000000000;
          rom[20] = 32'b00000000110111100100001010100000; // slt $9, $3, $7
          rom[21] = 32'b00000000001001100100000000000000;
          rom[22] = 32'b00101010011001000000000000000000; // slti $9, $0, -1 
          rom[23] = 32'b00000000001001100100000000000000;
          rom[24] = 32'b00001100001101000000000000000000; // jal 56
          rom[25] = 32'b00000000001101110100000000000000;
          rom[26] = 32'b00001000010011000000000000000000; // j 80
          rom[27] = 32'b00000000000011001100000000000000;
          rom[28] = 32'b01100000000001000000000001111100; // li $1, 31
          rom[29] = 32'b00000000000001000100000000000000;
          rom[30] = 32'b01100000000001000000000011111100; // li $1, 63
          rom[31] = 32'b00000000000001000100000000000000;
			 rom[32] = 32'b00000000100011000100001001010000; // or $1, $2, $3
          rom[33] = 32'b00000000000001000100000000000000;
          rom[34] = 32'b00000000100011000100001001000000; // and $1, $2, $3
          rom[35] = 32'b00000000000001000100000000000000; 
          rom[36] = 32'b00110000100001000000000000000100; // andi $1, $2, 1
          rom[37] = 32'b00000000000001000100000000000000;
			 rom[38] = 32'b00000000000111000101000000000000; // sll $1, $7, 4
          rom[39] = 32'b00000000000001000100000000000000;
          rom[40] = 32'b00110100100001000000000000010000; // ori $1, $2, 4
          rom[41] = 32'b00000000000001000100000000000000;
          rom[42] = 32'b00000000000101000100100000100000; // srl $1, $5, 2
          rom[43] = 32'b00000000000001000100000000000000;
			 rom[44] = 32'b00010110000000111111111111110100; // bne $8, $0, -3
          rom[45] = 32'b00000000000000000011110000000000;
          rom[46] = 32'b00010010000000000000000000000100; // beq $8, $0, 1
          rom[47] = 32'b00000000000000000000000000000000;
      end   
      assign instruction = rom[pc[10:1]];  
 endmodule 